module Registerfile(
    input [2:0] in,
    output []
);

endmodule