module filter(
    input [7:0]in1,
    input [7:0]in2,
    input [7:0]in3,
    input [7:0]in4,
    input [7:0]in5,
    input [7:0]in6,
    input [7:0]in7,
    input [7:0]in8,
    input ind,
    output reg [7:0] o1,
    output reg [7:0] o2,
    output reg [7:0] o3,
    output reg [7:0] o4,
    output reg [7:0] o5,
    output reg [7:0] o6,
    output reg [7:0] o7,
    output reg [7:0] o8
);
    

endmodule